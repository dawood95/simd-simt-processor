/*
 * Sheik Dawood
 * dawood0@purdue.edu
 * 
 * Vector load store unit
 */
